module alu
(
   	 input      [31:0] rs, rt, 
	 input	    [4:0] shamt, 
	 input	    [5:0] funct,
   	 output     [31:0] rd
);

	...
	
endmodule
